`include "1-IF_stage/InstructionRAM.v"

module IF_stage (
    input CLK

);
    
endmodule