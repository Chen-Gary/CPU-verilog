`include "InstructionRAM.v"

module IF_stage (
    input CLK,
    
);
    
endmodule